module hello_world();

	initial begin
	$display("\n\t hello world! \n");
	end

endmodule